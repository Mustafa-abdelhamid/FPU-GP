module Top_Add_Sub (

input     wire   [7:0]        Ex,Ey,
input     wire   [22:0]       Mx,My,
input     wire                Sx,Sy,EOP,sub,
input	  wire	 [1:0] 		  roundMode , ////
output    wire   [7:0]        Ez,
output    wire   [22:0]       Mz_final,
output    wire                Sz,
output	  wire  invalid_flag,overflow_flag,underflow_flag,inexact_flag,zero_flag ////////
); 
//////// LZA BLOCK  outputs ///////////
wire [26:0]E;
wire [4:0]SHL; // required left shift (may be wrong)
wire [26:0]sum_shifted;
wire second_shift_left;

wire [22:0]correct_sum_shifted;  //
//////// Exponent difference outputs ///////////
wire        sgn_d;
wire        zero_d;
wire [7:0]  d;

//////// Alignment outputs ///////////
wire [26:0] out_11;
wire [26:0] out_22;
wire  	    cmp;
//////// max exponent  outputs ///////////

wire [7:0]  maxOf_Ex_Ey;
//////// Exponent_Update  outputs ///////////
wire [4:0] mantissaReqiredModify ; // to modify mantisa in case of underflow
wire [7:0] Ez_updated;
wire overflow_case ; 
//underflow_flag  is output
//////// Mantissa MUX BLOCK  outputs /////////// 

wire [22:0]Mz_to_exceptions ;

wire       ovf;
wire  [4:0]final_shift_left;
wire ovf_rnd ;
/////////////////////////////////////////////////////////////////////////
////////////////////////////Exponent difference /////////////////////////
/////////////////////////////////////////////////////////////////////////



Exponent_Difference Ex_Diff (
.Ex(Ex),
.Ey(Ey),
.sgn_d(sgn_d),
.zero_d(zero_d),
.d(d)
);
////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////
////////////////////////////////Alignment  //////////////////////////////
/////////////////////////////////////////////////////////////////////////

Alignment A1 (
.Mx(Mx),
.My(My),
.sgn_d(sgn_d), 
.EOP(EOP),
.zero_d(zero_d),
.Ex(Ex),
.Ey(Ey),
.d(d),
.out_11(out_11),
.out_22(out_22),
.Cmp(cmp)
);

////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////
/////////////////////////////max exponent Mux  //////////////////////////
/////////////////////////////////////////////////////////////////////////


Mux mux11 (
.Ex(Ex),
.Ey(Ey),
.sgn_d(sgn_d),
.Out_mux(maxOf_Ex_Ey)
);
/////////////////////////////////////////////////////////////////////////


/////////////////////////////////////////////////////////////////////////
///////////////////////////// Exponent_Update  //////////////////////////
/////////////////////////////////////////////////////////////////////////

  

Exponent_Update Ex_update(
 .maxOf_Ex_Ey(maxOf_Ex_Ey), 
 .ovf(ovf),
 .ovf_rnd(ovf_rnd),///
 .reqiredShift_left(SHL) , // LZA output (shift requred for massive shifter)
 
 .mantissaReqiredModify (mantissaReqiredModify) , // to modify mantisa in case of underflow
 .Ez(Ez_updated),
 .underflow_flag(underflow_flag),
 .overflow_case(overflow_case) 
 );

//////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////
/////////////////////////////SIGN BLOCK  //////////////////////////
/////////////////////////////////////////////////////////////////////////

//////// SIGN BLOCK  outputs ///////////
//Sz is output 
Sign_of_z sign_z11 (
.Sx(Sx),
.Sy(Sy),
.EOP(EOP),
.cmp(cmp),
.sign_d(sgn_d),
.zero_d(zero_d),
.Sz(Sz)
);
//////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////
/////////////////////////////exceptions BLOCK  //////////////////////////
/////////////////////////////////////////////////////////////////////////

//////// exceptions BLOCK  outputs ///////////
// flags are outputs 
exceptions exceptions_block
 (.Ex (Ex),
 .Ey(Ey),
 .Mx(Mx),
 .My(My),
 .Mz(Mz_to_exceptions), /////Mn mantissa mux 
 .EOP(EOP),
 .exponent_z(Ez_updated),
 .overflow_case(overflow_case),
 
 .invalid_flag(invalid_flag),
 .overflow_flag(overflow_flag),
 .zero_flag(zero_flag)
 );
 
//////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////
/////////////////////////////adder BLOCK  //////////////////////////
/////////////////////////////////////////////////////////////////////////

//////// adder BLOCK  outputs ///////////
wire [26:0]sum;

wire [2:0] most_bits_of_adder_out ; 
 
adder_modified adder_mod_inst 
(
.A(out_11),
.B(out_22),
.sub(sub),
.sum(sum),
.ovf_out(ovf),
.most_bits_of_adder_out(most_bits_of_adder_out)
);

//////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////
/////////////////////////////LZA BLOCK  //////////////////////////
/////////////////////////////////////////////////////////////////////////



// // 
 
LZA_1_modified LZA_1_modified_inst (
.A(out_11),
.B(out_22),
.E(E)
);
  // generate E signal
LZA_2_modified LZA_2_modified_inst (
.E({ovf,E}),
.SHL(SHL)
); // count number of Zeros

first_massive_shift_left first_massive_shift_left_inst (
.adder_out(sum) , 
.SHL(SHL) , 
.sum_shifted( sum_shifted)
);  // shift sum by the required amount
 
LZA_final_modified LZA_final_modified_inst ( 
.sum_shifted(sum_shifted) ,
.correct_sum_shifted (correct_sum_shifted) , 
.second_shift_left (second_shift_left)

 ); // check for correctness 
 

shift_left_adder shift_left_adder_inst (
.SHL(SHL) ,
.second_shift_left(second_shift_left) , 
.final_shift_left(final_shift_left)

 ); //modify in case of error 

/////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////
//////////////////////// L1/R1 shifter BLOCK  ///////////////////////////
/////////////////////////////////////////////////////////////////////////

//////// L1/R1 shifter BLOCK  outputs ///////////
wire [26:0]righPass_shift_out;  
wire [1:0]righPath_exponentUpdate_control;

left_right_shifter left_right_shifter_inst (
.adder_out(sum) , 
.ovf(ovf) , 
.righPass_shift_out(righPass_shift_out),
.righPath_exponentUpdate_control (righPath_exponentUpdate_control) 

 );

/////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////
//////////////////////// ROUND BLOCK  ///////////////////////////
/////////////////////////////////////////////////////////////////////////

//////// ROUND BLOCK  outputs ///////////
wire [22:0] rounded_mantissa;
// 
// inexact flag is output 
ROUND ROUND_inst ( 
.Min(righPass_shift_out)   ,
.roundMode (roundMode),		
.Sign_in(Sz) ,

.MOut (rounded_mantissa)  ,
.overFlow(ovf_rnd),
.inexact_flag(inexact_flag)
);

/////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////
//////////////////////// Mantissa MUX BLOCK  ///////////////////////////
/////////////////////////////////////////////////////////////////////////


 
mantessa_mux mantessa_mux_inst (
.left_path (correct_sum_shifted),
.right_path (rounded_mantissa) , 
.most_bits_of_adder_out(most_bits_of_adder_out) , 
.final_mantessa (Mz_to_exceptions)
 );
 
 
final_output final_output_inst (
.M_out (Mz_to_exceptions) ,
.E_out(Ez_updated) ,
.required_modify (final_shift_left)  ,

.overflow_flag(overflow_flag) , 
.underflow_flag(underflow_flag) , 
.invalid_flag(invalid_flag) , 

.final_M_out (Mz_final) ,
.final_E_out (Ez)

);
 
 
 endmodule
