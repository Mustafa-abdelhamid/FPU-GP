module normalization 

(
input 	wire				CLK,RST,
input	wire	[47:0]		P,
input	wire	[9:0] 		Ez_add,
output	reg 	[24:0]		normalised_output , // hidden + 23 mantissa + sticky bit 
output 	reg 	[4:0] 		SHL ,
output 	reg 				ovf  ,
output	reg		[46:0] 		after_sh_norm
);

wire	 [9:0] 		den_exponent    ; 
wire				handel_464_case ;

reg	[47:0]		P_ff;

reg	[9:0] 		EzAdd_f,EzAdd_ff;



assign handel_464_case = ~|EzAdd_ff    ;
assign den_exponent = ~EzAdd_ff + 1'b1 ;


always @ (posedge CLK or negedge RST )
	begin
	if (!RST) 
		begin
////////inputs RST
			P_ff 		<= 0;
			EzAdd_f		<= 0;
			EzAdd_ff	<= 0;
		end
		
	else
		begin
////////inputs Reg
			P_ff 		<= P ;
			EzAdd_f		<= Ez_add ;
			EzAdd_ff	<= EzAdd_f ;

		end			
	end


always@(*)

begin 
	if (!EzAdd_ff[9] & !handel_464_case)
	begin
	if (!P_ff[47])  // already normalised or Leading zeros
		begin
		ovf = 1'b0 ;
		casez(P_ff[46:0]) // synopsys full_case parallel_case
				47'b1?????????????????????????????????????????????? : // already normalised
					begin
						SHL = 0;
						after_sh_norm = P_ff[46:0];
						normalised_output= after_sh_norm[46:22] ; 
					end
				47'b01????????????????????????????????????????????? : // leading zero 
					begin
						SHL = 1;
						after_sh_norm = P_ff[46:0]<<1;
						normalised_output= after_sh_norm[46:22] ; 
					end
				
				47'b001???????????????????????????????????????????? : // leading zero 
					begin
						SHL = 2;
						after_sh_norm = P_ff[46:0]<<2;
						normalised_output= after_sh_norm[46:22] ; 
					end
				
				47'b0001??????????????????????????????????????????? : // leading zero 
					begin
						SHL = 3;
						after_sh_norm = P_ff[46:0]<<3;
						normalised_output= after_sh_norm[46:22] ; 
					end
				
				47'b00001?????????????????????????????????????????? : // leading zero 
					begin
						SHL = 4;
						after_sh_norm = P_ff[46:0]<<4;
						normalised_output= after_sh_norm[46:22] ;  
					end
					
				47'b000001????????????????????????????????????????? : // leading zero
					begin
						SHL = 5;
						after_sh_norm = P_ff[46:0]<<5;
						normalised_output= after_sh_norm[46:22] ;  
					end
				
				47'b0000001???????????????????????????????????????? : // leading zero
					begin
						SHL = 6;
						after_sh_norm = P_ff[46:0]<<6;
						normalised_output= after_sh_norm[46:22] ; 
					end
				47'b00000001??????????????????????????????????????? : // leading zero
					begin
						SHL = 7;
						after_sh_norm = P_ff[46:0]<<7;
						normalised_output= after_sh_norm[46:22] ; 
					end
				47'b000000001?????????????????????????????????????? : // leading zero
					begin
						SHL = 8;
						after_sh_norm = P_ff[46:0]<<8;
						normalised_output= after_sh_norm[46:22] ; 
					end
				47'b0000000001????????????????????????????????????? : // leading zero
					begin
						SHL = 9;
						after_sh_norm = P_ff[46:0]<<9;
						normalised_output= after_sh_norm[46:22] ; 
					end
				47'b00000000001???????????????????????????????????? : // leading zero
					begin
						SHL = 10;
						after_sh_norm = P_ff[46:0]<<10;
						normalised_output= after_sh_norm[46:22] ;  
					end
				47'b0000_0000_0001_????_????_????_??????????????????????? : // leading zero
					begin
						SHL = 11;
						after_sh_norm = P_ff[46:0]<<11;
						normalised_output= after_sh_norm[46:22] ; 
					end
				
				47'b0000_0000_0000_1???_????_????_??????????????????????? : // leading zero
					begin
						SHL = 12;
						after_sh_norm = P_ff[46:0]<<12;
						normalised_output= after_sh_norm[46:22] ; 
					end
				
				47'b0000_0000_0000_01??_????_????_??????????????????????? : // leading zero
					begin
						SHL = 13;
						after_sh_norm = P_ff[46:0]<<13;
						normalised_output= after_sh_norm[46:22] ; 
					end
				
				47'b0000_0000_0000_001?_????_????_??????????????????????? : // leading zero
					begin
						SHL = 14;
						after_sh_norm = P_ff[46:0]<<14;
						normalised_output= after_sh_norm[46:22] ;  
					end
				
				47'b0000_0000_0000_0001_????_????_??????????????????????? : // leading zero
					begin
						SHL = 15;
						after_sh_norm = P_ff[46:0]<<15;
						normalised_output= after_sh_norm[46:22] ; 
					end
				
				47'b0000_0000_0000_0000_1???_????_??????????????????????? : // leading zero
					begin
						SHL = 16;
						after_sh_norm = P_ff[46:0]<<16;
						normalised_output= after_sh_norm[46:22] ;  
					end
				
				47'b0000_0000_0000_0000_01??_????_??????????????????????? : // leading zero
					begin
						SHL = 17;
						after_sh_norm = P_ff[46:0]<<17;
						normalised_output= after_sh_norm[46:22] ; 
					end
				
				47'b0000_0000_0000_0000_001?_????_??????????????????????? : // leading zero
					begin
						SHL = 18;
						after_sh_norm = P_ff[46:0]<<18;
						normalised_output= after_sh_norm[46:22] ; 
					end
				
								
				47'b0000_0000_0000_0000_0001_????_??????????????????????? : // leading zero
					begin
						SHL = 19;
						after_sh_norm = P_ff[46:0]<<19;
						normalised_output= after_sh_norm[46:22] ; 
					end
								
				47'b0000_0000_0000_0000_0000_1???_??????????????????????? : // leading zero
					begin
						SHL = 20;
						after_sh_norm = P_ff[46:0]<<20;
						normalised_output= after_sh_norm[46:22] ; 
					end
				
								
				47'b0000_0000_0000_0000_0000_01??_??????????????????????? : // leading zero
					begin
						SHL = 21;
						after_sh_norm = P_ff[46:0]<<21;
						normalised_output= after_sh_norm[46:22] ; 
					end
								
				47'b0000_0000_0000_0000_0000_001?_??????????????????????? : // leading zero
					begin
						SHL = 22;
						after_sh_norm = P_ff[46:0]<<22;
						normalised_output= after_sh_norm[46:22] ; 
					end
				
				47'b0000_0000_0000_0000_0000_0001_??????????????????????? : // leading zero
					begin
						SHL = 23;
						after_sh_norm = P_ff[46:0]<<23;
						normalised_output= after_sh_norm[46:22] ;  
					end
				47'b0000_0000_0000_0000_0000_0000_1?????????????????????? : // leading zero
					begin
						SHL = 24;
						after_sh_norm = P_ff[46:0]<<24;
						normalised_output= after_sh_norm[46:22] ; 
					end
				
				endcase
		  
		end 
	else 
		begin
			SHL=0 ;
			ovf= 1'b1 ;
			after_sh_norm = P_ff[46:0];
			normalised_output= P_ff [47:23] ; 
		end 
	end
	
	else  /// incase of negative exponent
		begin
				SHL=0 ;
				after_sh_norm = P_ff[47:1]; //// very important range ?????????????????
				ovf= P_ff[47] ;
				normalised_output = P_ff [47:23] >> den_exponent ;

		end
end 

endmodule